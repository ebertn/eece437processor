`include "forward_if.vh"
`include "cpu_types_pkg.vh"

module forward_unit
(
	forward_if forif
); 


import cpu_types_pkg::*;



endmodule
