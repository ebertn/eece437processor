module ex_mem
(

); 