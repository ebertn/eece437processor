

module if_id 
(
	


); 