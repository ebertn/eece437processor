module mem_wb
(

); 