module id_ex
(

); 
