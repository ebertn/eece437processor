`include "cpu_types_pkg.vh"
`include "register_file_if.vh"

module register_file (
  input logic CLK,
  nRST,
  register_file_if.rf rfif
);

import cpu_types_pkg::*;

word_t [31:0] registers, next_registers;

always_ff @(posedge CLK, negedge nRST) begin
	if (!nRST) begin
		registers <= '0;
	end else begin
		registers <= next_registers;
	end
end

always_comb begin
	//next_registers = '0;

	next_registers = registers;
	next_registers[rfif.wsel] = rfif.WEN ? rfif.wdat : registers[rfif.wsel];
	next_registers[0] = '0;

	rfif.rdat1 = registers[rfif.rsel1];
	rfif.rdat2 = registers[rfif.rsel2];
end

endmodule